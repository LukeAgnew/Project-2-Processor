library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity memory_m_16bit is
    Port ( address : in  unsigned STD_LOGIC_VECTOR (15 downto 0);
           write_data : in  STD_LOGIC_VECTOR (15 downto 0);
           MemWrite, MemRead : in  STD_LOGIC;
			  Clk : in STD_LOGIC;
           read_data : out  STD_LOGIC_VECTOR (15 downto 0));
end memory_m_16bit;

architecture Behavioral of memory_m_16bit is
type mem_array is array(0 to 511) of std_logic_vector(15 downto 0);
-- define type, for memory arrays
begin
	mem_process: process (address, write_data)
	-- initialize data memory, X denotes hexadecimal number
	variable data_mem : mem_array := (
			-- 0
			X"0000", -- 0 
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7

			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
			
			-- 1
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
				
			-- 2
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 3
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 4
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 5
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 6
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 7
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 8
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 9
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
			
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- A
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- B
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
				
			-- C
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- D
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
			
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
				
			-- E
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- F
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
			
			
			-- 10
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
			
			-- 11
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
			-- 12
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
			
			-- 13
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 14
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
			
			-- 15
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
		
			-- 16
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 17
		X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
			
			-- 18
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 19
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
			
			-- 1A
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 1B
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
			
			-- 1C
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
		
			-- 1D
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F
			
			-- 1E
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000", -- F

			-- 1F
			X"0000", -- 0
			X"0000", -- 1
			X"0000", -- 2
			X"0000", -- 3
			X"0000", -- 4
			X"0000", -- 5
			X"0000", -- 6
			X"0000", -- 7
				
			X"0000", -- 8
			X"0000", -- 9
			X"0000", -- A
			X"0000", -- B
			X"0000", -- C
			X"0000", -- D
			X"0000", -- E
			X"0000" -- F
			);
	variable addr:integer;
	begin -- the following type conversion function is in std_logic_arith
		addr:=conv_integer(address(2 downto 0));
		if MemWrite ='1' then
			data_mem(addr):= write_data;
		elsif MemRead='1' then
			read_data <= data_mem(addr) after 10 ns;
		end if;
	end process;

end Behavioral;

